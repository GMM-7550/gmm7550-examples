
library ieee;
use ieee.std_logic_1164.all;

package bcm_pkg is
  type std_logic_vector_array_t is array (natural range <>) of std_logic_vector;
end package bcm_pkg;
