../../blink_25/src/blink.vhd